library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ide_cffa_rom is
port (
	clk  : in  std_logic;
	addr : in  unsigned(11 downto 0);
	data : out unsigned(7 downto 0)
);
end entity;

architecture prom of ide_cffa_rom is
	type rom is array(0 to  4095) of unsigned(7 downto 0);
	signal rom_data: rom := (
		X"43",X"46",X"46",X"41",X"20",X"46",X"69",X"72",X"6D",X"77",X"61",X"72",X"65",X"0D",X"0D",X"0D",
		X"53",X"65",X"65",X"20",X"3C",X"68",X"74",X"74",X"70",X"3A",X"2F",X"2F",X"64",X"72",X"65",X"68",
		X"65",X"72",X"2E",X"6E",X"65",X"74",X"2F",X"43",X"46",X"66",X"6F",X"72",X"41",X"70",X"70",X"6C",
		X"65",X"49",X"49",X"2F",X"3E",X"2E",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",
		X"56",X"65",X"72",X"73",X"69",X"6F",X"6E",X"20",X"32",X"2E",X"30",X"20",X"66",X"6F",X"72",X"20",
		X"36",X"35",X"30",X"32",X"20",X"6F",X"72",X"20",X"6C",X"61",X"74",X"65",X"72",X"2E",X"0D",X"0D",
		X"52",X"65",X"71",X"75",X"69",X"72",X"65",X"73",X"20",X"43",X"46",X"46",X"41",X"20",X"77",X"69",
		X"74",X"68",X"20",X"45",X"45",X"50",X"52",X"4F",X"4D",X"2C",X"20",X"6E",X"6F",X"74",X"20",X"45",
		X"50",X"52",X"4F",X"4D",X"2E",X"0D",X"0D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"A9",X"20",X"A2",X"00",X"A9",X"03",X"A9",X"3C",X"10",X"0A",X"18",X"90",X"01",X"38",X"20",X"A1",
		X"C1",X"4C",X"28",X"C8",X"20",X"A1",X"C1",X"86",X"43",X"AC",X"0B",X"C8",X"A9",X"C5",X"20",X"A8",
		X"FC",X"88",X"D0",X"F8",X"AD",X"00",X"C0",X"2D",X"09",X"C8",X"CD",X"0A",X"C8",X"D0",X"07",X"EA",
		X"20",X"A1",X"C1",X"20",X"2B",X"C8",X"A0",X"01",X"84",X"42",X"88",X"84",X"46",X"84",X"47",X"A9",
		X"08",X"85",X"45",X"84",X"44",X"20",X"A1",X"C1",X"20",X"37",X"C8",X"85",X"FF",X"B0",X"10",X"AC",
		X"00",X"08",X"88",X"D0",X"0A",X"AD",X"01",X"08",X"F0",X"05",X"A6",X"43",X"4C",X"01",X"08",X"A5",
		X"00",X"D0",X"0A",X"A5",X"01",X"CD",X"F8",X"07",X"D0",X"03",X"4C",X"BA",X"FA",X"20",X"2E",X"C8",
		X"A0",X"00",X"A6",X"FF",X"D0",X"02",X"A0",X"0E",X"20",X"95",X"C1",X"8A",X"F0",X"0C",X"AD",X"79",
		X"07",X"0A",X"0A",X"A9",X"B0",X"69",X"00",X"20",X"ED",X"FD",X"A0",X"1C",X"20",X"95",X"C1",X"20",
		X"A1",X"C1",X"4C",X"34",X"C8",X"B9",X"BC",X"C1",X"F0",X"06",X"20",X"31",X"C8",X"C8",X"D0",X"F5",
		X"60",X"8D",X"92",X"C0",X"A9",X"C1",X"8D",X"F8",X"07",X"2C",X"FF",X"CF",X"AD",X"20",X"C8",X"49",
		X"CF",X"D0",X"05",X"A0",X"01",X"A2",X"10",X"60",X"20",X"93",X"FE",X"00",X"43",X"68",X"65",X"63",
		X"6B",X"20",X"64",X"65",X"76",X"69",X"63",X"65",X"20",X"00",X"4E",X"6F",X"20",X"62",X"6F",X"6F",
		X"74",X"20",X"62",X"6C",X"6F",X"63",X"6B",X"00",X"2E",X"0D",X"0D",X"43",X"6F",X"75",X"6C",X"64",
		X"20",X"6E",X"6F",X"74",X"20",X"62",X"6F",X"6F",X"74",X"20",X"70",X"61",X"72",X"74",X"69",X"74",
		X"69",X"6F",X"6E",X"20",X"00",X"FF",X"43",X"46",X"46",X"41",X"FF",X"00",X"00",X"00",X"17",X"0A",
		X"A9",X"20",X"A2",X"00",X"A9",X"03",X"A9",X"3C",X"10",X"0A",X"18",X"90",X"01",X"38",X"20",X"A1",
		X"C2",X"4C",X"28",X"C8",X"20",X"A1",X"C2",X"86",X"43",X"AC",X"0B",X"C8",X"A9",X"C5",X"20",X"A8",
		X"FC",X"88",X"D0",X"F8",X"AD",X"00",X"C0",X"2D",X"09",X"C8",X"CD",X"0A",X"C8",X"D0",X"07",X"EA",
		X"20",X"A1",X"C2",X"20",X"2B",X"C8",X"A0",X"01",X"84",X"42",X"88",X"84",X"46",X"84",X"47",X"A9",
		X"08",X"85",X"45",X"84",X"44",X"20",X"A1",X"C2",X"20",X"37",X"C8",X"85",X"FF",X"B0",X"10",X"AC",
		X"00",X"08",X"88",X"D0",X"0A",X"AD",X"01",X"08",X"F0",X"05",X"A6",X"43",X"4C",X"01",X"08",X"A5",
		X"00",X"D0",X"0A",X"A5",X"01",X"CD",X"F8",X"07",X"D0",X"03",X"4C",X"BA",X"FA",X"20",X"2E",X"C8",
		X"A0",X"00",X"A6",X"FF",X"D0",X"02",X"A0",X"0E",X"20",X"95",X"C2",X"8A",X"F0",X"0C",X"AD",X"7A",
		X"07",X"0A",X"0A",X"A9",X"B0",X"69",X"00",X"20",X"ED",X"FD",X"A0",X"1C",X"20",X"95",X"C2",X"20",
		X"A1",X"C2",X"4C",X"34",X"C8",X"B9",X"BC",X"C2",X"F0",X"06",X"20",X"31",X"C8",X"C8",X"D0",X"F5",
		X"60",X"8D",X"A2",X"C0",X"A9",X"C2",X"8D",X"F8",X"07",X"2C",X"FF",X"CF",X"AD",X"20",X"C8",X"49",
		X"CF",X"D0",X"05",X"A0",X"02",X"A2",X"20",X"60",X"20",X"93",X"FE",X"00",X"43",X"68",X"65",X"63",
		X"6B",X"20",X"64",X"65",X"76",X"69",X"63",X"65",X"20",X"00",X"4E",X"6F",X"20",X"62",X"6F",X"6F",
		X"74",X"20",X"62",X"6C",X"6F",X"63",X"6B",X"00",X"2E",X"0D",X"0D",X"43",X"6F",X"75",X"6C",X"64",
		X"20",X"6E",X"6F",X"74",X"20",X"62",X"6F",X"6F",X"74",X"20",X"70",X"61",X"72",X"74",X"69",X"74",
		X"69",X"6F",X"6E",X"20",X"00",X"FF",X"43",X"46",X"46",X"41",X"FF",X"00",X"00",X"00",X"17",X"0A",
		X"A9",X"20",X"A2",X"00",X"A9",X"03",X"A9",X"3C",X"10",X"0A",X"18",X"90",X"01",X"38",X"20",X"A1",
		X"C3",X"4C",X"28",X"C8",X"20",X"A1",X"C3",X"86",X"43",X"AC",X"0B",X"C8",X"A9",X"C5",X"20",X"A8",
		X"FC",X"88",X"D0",X"F8",X"AD",X"00",X"C0",X"2D",X"09",X"C8",X"CD",X"0A",X"C8",X"D0",X"07",X"EA",
		X"20",X"A1",X"C3",X"20",X"2B",X"C8",X"A0",X"01",X"84",X"42",X"88",X"84",X"46",X"84",X"47",X"A9",
		X"08",X"85",X"45",X"84",X"44",X"20",X"A1",X"C3",X"20",X"37",X"C8",X"85",X"FF",X"B0",X"10",X"AC",
		X"00",X"08",X"88",X"D0",X"0A",X"AD",X"01",X"08",X"F0",X"05",X"A6",X"43",X"4C",X"01",X"08",X"A5",
		X"00",X"D0",X"0A",X"A5",X"01",X"CD",X"F8",X"07",X"D0",X"03",X"4C",X"BA",X"FA",X"20",X"2E",X"C8",
		X"A0",X"00",X"A6",X"FF",X"D0",X"02",X"A0",X"0E",X"20",X"95",X"C3",X"8A",X"F0",X"0C",X"AD",X"7B",
		X"07",X"0A",X"0A",X"A9",X"B0",X"69",X"00",X"20",X"ED",X"FD",X"A0",X"1C",X"20",X"95",X"C3",X"20",
		X"A1",X"C3",X"4C",X"34",X"C8",X"B9",X"BC",X"C3",X"F0",X"06",X"20",X"31",X"C8",X"C8",X"D0",X"F5",
		X"60",X"8D",X"B2",X"C0",X"A9",X"C3",X"8D",X"F8",X"07",X"2C",X"FF",X"CF",X"AD",X"20",X"C8",X"49",
		X"CF",X"D0",X"05",X"A0",X"03",X"A2",X"30",X"60",X"20",X"93",X"FE",X"00",X"43",X"68",X"65",X"63",
		X"6B",X"20",X"64",X"65",X"76",X"69",X"63",X"65",X"20",X"00",X"4E",X"6F",X"20",X"62",X"6F",X"6F",
		X"74",X"20",X"62",X"6C",X"6F",X"63",X"6B",X"00",X"2E",X"0D",X"0D",X"43",X"6F",X"75",X"6C",X"64",
		X"20",X"6E",X"6F",X"74",X"20",X"62",X"6F",X"6F",X"74",X"20",X"70",X"61",X"72",X"74",X"69",X"74",
		X"69",X"6F",X"6E",X"20",X"00",X"FF",X"43",X"46",X"46",X"41",X"FF",X"00",X"00",X"00",X"17",X"0A",
		X"A9",X"20",X"A2",X"00",X"A9",X"03",X"A9",X"3C",X"10",X"0A",X"18",X"90",X"01",X"38",X"20",X"A1",
		X"C4",X"4C",X"28",X"C8",X"20",X"A1",X"C4",X"86",X"43",X"AC",X"0B",X"C8",X"A9",X"C5",X"20",X"A8",
		X"FC",X"88",X"D0",X"F8",X"AD",X"00",X"C0",X"2D",X"09",X"C8",X"CD",X"0A",X"C8",X"D0",X"07",X"EA",
		X"20",X"A1",X"C4",X"20",X"2B",X"C8",X"A0",X"01",X"84",X"42",X"88",X"84",X"46",X"84",X"47",X"A9",
		X"08",X"85",X"45",X"84",X"44",X"20",X"A1",X"C4",X"20",X"37",X"C8",X"85",X"FF",X"B0",X"10",X"AC",
		X"00",X"08",X"88",X"D0",X"0A",X"AD",X"01",X"08",X"F0",X"05",X"A6",X"43",X"4C",X"01",X"08",X"A5",
		X"00",X"D0",X"0A",X"A5",X"01",X"CD",X"F8",X"07",X"D0",X"03",X"4C",X"BA",X"FA",X"20",X"2E",X"C8",
		X"A0",X"00",X"A6",X"FF",X"D0",X"02",X"A0",X"0E",X"20",X"95",X"C4",X"8A",X"F0",X"0C",X"AD",X"7C",
		X"07",X"0A",X"0A",X"A9",X"B0",X"69",X"00",X"20",X"ED",X"FD",X"A0",X"1C",X"20",X"95",X"C4",X"20",
		X"A1",X"C4",X"4C",X"34",X"C8",X"B9",X"BC",X"C4",X"F0",X"06",X"20",X"31",X"C8",X"C8",X"D0",X"F5",
		X"60",X"8D",X"C2",X"C0",X"A9",X"C4",X"8D",X"F8",X"07",X"2C",X"FF",X"CF",X"AD",X"20",X"C8",X"49",
		X"CF",X"D0",X"05",X"A0",X"04",X"A2",X"40",X"60",X"20",X"93",X"FE",X"00",X"43",X"68",X"65",X"63",
		X"6B",X"20",X"64",X"65",X"76",X"69",X"63",X"65",X"20",X"00",X"4E",X"6F",X"20",X"62",X"6F",X"6F",
		X"74",X"20",X"62",X"6C",X"6F",X"63",X"6B",X"00",X"2E",X"0D",X"0D",X"43",X"6F",X"75",X"6C",X"64",
		X"20",X"6E",X"6F",X"74",X"20",X"62",X"6F",X"6F",X"74",X"20",X"70",X"61",X"72",X"74",X"69",X"74",
		X"69",X"6F",X"6E",X"20",X"00",X"FF",X"43",X"46",X"46",X"41",X"FF",X"00",X"00",X"00",X"17",X"0A",
		X"A9",X"20",X"A2",X"00",X"A9",X"03",X"A9",X"00",X"10",X"0A",X"18",X"90",X"01",X"38",X"20",X"A1",
		X"C5",X"4C",X"28",X"C8",X"20",X"A1",X"C5",X"86",X"43",X"AC",X"0B",X"C8",X"A9",X"C5",X"20",X"A8",
		X"FC",X"88",X"D0",X"F8",X"AD",X"00",X"C0",X"2D",X"09",X"C8",X"CD",X"0A",X"C8",X"D0",X"07",X"EA",
		X"20",X"A1",X"C5",X"20",X"2B",X"C8",X"A0",X"01",X"84",X"42",X"88",X"84",X"46",X"84",X"47",X"A9",
		X"08",X"85",X"45",X"84",X"44",X"20",X"A1",X"C5",X"20",X"37",X"C8",X"85",X"FF",X"B0",X"10",X"AC",
		X"00",X"08",X"88",X"D0",X"0A",X"AD",X"01",X"08",X"F0",X"05",X"A6",X"43",X"4C",X"01",X"08",X"A5",
		X"00",X"D0",X"0A",X"A5",X"01",X"CD",X"F8",X"07",X"D0",X"03",X"4C",X"BA",X"FA",X"20",X"2E",X"C8",
		X"A0",X"00",X"A6",X"FF",X"D0",X"02",X"A0",X"0E",X"20",X"95",X"C5",X"8A",X"F0",X"0C",X"AD",X"7D",
		X"07",X"0A",X"0A",X"A9",X"B0",X"69",X"00",X"20",X"ED",X"FD",X"A0",X"1C",X"20",X"95",X"C5",X"20",
		X"A1",X"C5",X"4C",X"34",X"C8",X"B9",X"BC",X"C5",X"F0",X"06",X"20",X"31",X"C8",X"C8",X"D0",X"F5",
		X"60",X"8D",X"D2",X"C0",X"A9",X"C5",X"8D",X"F8",X"07",X"2C",X"FF",X"CF",X"AD",X"20",X"C8",X"49",
		X"CF",X"D0",X"05",X"A0",X"05",X"A2",X"50",X"60",X"20",X"93",X"FE",X"00",X"43",X"68",X"65",X"63",
		X"6B",X"20",X"64",X"65",X"76",X"69",X"63",X"65",X"20",X"00",X"4E",X"6F",X"20",X"62",X"6F",X"6F",
		X"74",X"20",X"62",X"6C",X"6F",X"63",X"6B",X"00",X"2E",X"0D",X"0D",X"43",X"6F",X"75",X"6C",X"64",
		X"20",X"6E",X"6F",X"74",X"20",X"62",X"6F",X"6F",X"74",X"20",X"70",X"61",X"72",X"74",X"69",X"74",
		X"69",X"6F",X"6E",X"20",X"00",X"FF",X"43",X"46",X"46",X"41",X"FF",X"00",X"00",X"00",X"17",X"0A",
		X"A9",X"20",X"A2",X"00",X"A9",X"03",X"A9",X"3C",X"10",X"0A",X"18",X"90",X"01",X"38",X"20",X"A1",
		X"C6",X"4C",X"28",X"C8",X"20",X"A1",X"C6",X"86",X"43",X"AC",X"0B",X"C8",X"A9",X"C5",X"20",X"A8",
		X"FC",X"88",X"D0",X"F8",X"AD",X"00",X"C0",X"2D",X"09",X"C8",X"CD",X"0A",X"C8",X"D0",X"07",X"EA",
		X"20",X"A1",X"C6",X"20",X"2B",X"C8",X"A0",X"01",X"84",X"42",X"88",X"84",X"46",X"84",X"47",X"A9",
		X"08",X"85",X"45",X"84",X"44",X"20",X"A1",X"C6",X"20",X"37",X"C8",X"85",X"FF",X"B0",X"10",X"AC",
		X"00",X"08",X"88",X"D0",X"0A",X"AD",X"01",X"08",X"F0",X"05",X"A6",X"43",X"4C",X"01",X"08",X"A5",
		X"00",X"D0",X"0A",X"A5",X"01",X"CD",X"F8",X"07",X"D0",X"03",X"4C",X"BA",X"FA",X"20",X"2E",X"C8",
		X"A0",X"00",X"A6",X"FF",X"D0",X"02",X"A0",X"0E",X"20",X"95",X"C6",X"8A",X"F0",X"0C",X"AD",X"7E",
		X"07",X"0A",X"0A",X"A9",X"B0",X"69",X"00",X"20",X"ED",X"FD",X"A0",X"1C",X"20",X"95",X"C6",X"20",
		X"A1",X"C6",X"4C",X"34",X"C8",X"B9",X"BC",X"C6",X"F0",X"06",X"20",X"31",X"C8",X"C8",X"D0",X"F5",
		X"60",X"8D",X"E2",X"C0",X"A9",X"C6",X"8D",X"F8",X"07",X"2C",X"FF",X"CF",X"AD",X"20",X"C8",X"49",
		X"CF",X"D0",X"05",X"A0",X"06",X"A2",X"60",X"60",X"20",X"93",X"FE",X"00",X"43",X"68",X"65",X"63",
		X"6B",X"20",X"64",X"65",X"76",X"69",X"63",X"65",X"20",X"00",X"4E",X"6F",X"20",X"62",X"6F",X"6F",
		X"74",X"20",X"62",X"6C",X"6F",X"63",X"6B",X"00",X"2E",X"0D",X"0D",X"43",X"6F",X"75",X"6C",X"64",
		X"20",X"6E",X"6F",X"74",X"20",X"62",X"6F",X"6F",X"74",X"20",X"70",X"61",X"72",X"74",X"69",X"74",
		X"69",X"6F",X"6E",X"20",X"00",X"FF",X"43",X"46",X"46",X"41",X"FF",X"00",X"00",X"00",X"17",X"0A",
		X"A9",X"20",X"A2",X"00",X"A9",X"03",X"A9",X"3C",X"10",X"0A",X"18",X"90",X"01",X"38",X"20",X"A1",
		X"C7",X"4C",X"28",X"C8",X"20",X"A1",X"C7",X"86",X"43",X"AC",X"0B",X"C8",X"A9",X"C5",X"20",X"A8",
		X"FC",X"88",X"D0",X"F8",X"AD",X"00",X"C0",X"2D",X"09",X"C8",X"CD",X"0A",X"C8",X"D0",X"07",X"EA",
		X"20",X"A1",X"C7",X"20",X"2B",X"C8",X"A0",X"01",X"84",X"42",X"88",X"84",X"46",X"84",X"47",X"A9",
		X"08",X"85",X"45",X"84",X"44",X"20",X"A1",X"C7",X"20",X"37",X"C8",X"85",X"FF",X"B0",X"10",X"AC",
		X"00",X"08",X"88",X"D0",X"0A",X"AD",X"01",X"08",X"F0",X"05",X"A6",X"43",X"4C",X"01",X"08",X"A5",
		X"00",X"D0",X"0A",X"A5",X"01",X"CD",X"F8",X"07",X"D0",X"03",X"4C",X"BA",X"FA",X"20",X"2E",X"C8",
		X"A0",X"00",X"A6",X"FF",X"D0",X"02",X"A0",X"0E",X"20",X"95",X"C7",X"8A",X"F0",X"0C",X"AD",X"7F",
		X"07",X"0A",X"0A",X"A9",X"B0",X"69",X"00",X"20",X"ED",X"FD",X"A0",X"1C",X"20",X"95",X"C7",X"20",
		X"A1",X"C7",X"4C",X"34",X"C8",X"B9",X"BC",X"C7",X"F0",X"06",X"20",X"31",X"C8",X"C8",X"D0",X"F5",
		X"60",X"8D",X"F2",X"C0",X"A9",X"C7",X"8D",X"F8",X"07",X"2C",X"FF",X"CF",X"AD",X"20",X"C8",X"49",
		X"CF",X"D0",X"05",X"A0",X"07",X"A2",X"70",X"60",X"20",X"93",X"FE",X"00",X"43",X"68",X"65",X"63",
		X"6B",X"20",X"64",X"65",X"76",X"69",X"63",X"65",X"20",X"00",X"4E",X"6F",X"20",X"62",X"6F",X"6F",
		X"74",X"20",X"62",X"6C",X"6F",X"63",X"6B",X"00",X"2E",X"0D",X"0D",X"43",X"6F",X"75",X"6C",X"64",
		X"20",X"6E",X"6F",X"74",X"20",X"62",X"6F",X"6F",X"74",X"20",X"70",X"61",X"72",X"74",X"69",X"74",
		X"69",X"6F",X"6E",X"20",X"00",X"FF",X"43",X"46",X"46",X"41",X"FF",X"00",X"00",X"00",X"17",X"0A",
		X"04",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"DF",X"CD",X"05",X"1F",X"64",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"CF",X"FA",X"20",X"11",X"C0",X"00",X"00",X"07",X"4C",X"B9",X"CA",X"4C",X"1E",X"CE",X"4C",X"59",
		X"C8",X"4C",X"84",X"CF",X"4C",X"3A",X"C8",X"4C",X"BE",X"CA",X"B9",X"F8",X"07",X"18",X"69",X"01",
		X"20",X"6D",X"CF",X"20",X"8E",X"FD",X"20",X"DD",X"FB",X"A6",X"FF",X"F0",X"09",X"A0",X"15",X"20",
		X"61",X"CF",X"8A",X"20",X"DA",X"FD",X"4C",X"00",X"E0",X"20",X"2F",X"FB",X"20",X"84",X"FE",X"20",
		X"58",X"FC",X"20",X"93",X"FE",X"20",X"89",X"FE",X"20",X"81",X"C8",X"A0",X"00",X"20",X"61",X"CF",
		X"A9",X"22",X"85",X"24",X"A0",X"0E",X"20",X"61",X"CF",X"AD",X"F8",X"07",X"49",X"70",X"20",X"ED",
		X"FD",X"A0",X"28",X"A9",X"AD",X"20",X"ED",X"FD",X"88",X"D0",X"F8",X"60",X"A0",X"0C",X"B9",X"40",
		X"00",X"48",X"88",X"10",X"F9",X"86",X"41",X"BA",X"BD",X"0E",X"01",X"85",X"48",X"18",X"69",X"03",
		X"9D",X"0E",X"01",X"BD",X"0F",X"01",X"85",X"49",X"69",X"00",X"9D",X"0F",X"01",X"AD",X"F8",X"07",
		X"29",X"0F",X"85",X"40",X"A8",X"A6",X"41",X"20",X"FB",X"CB",X"A0",X"01",X"B1",X"48",X"85",X"42",
		X"C8",X"B1",X"48",X"AA",X"C8",X"B1",X"48",X"85",X"49",X"86",X"48",X"A9",X"01",X"A6",X"42",X"E0",
		X"0A",X"B0",X"1C",X"A0",X"00",X"B1",X"48",X"DD",X"10",X"C9",X"D0",X"27",X"A0",X"01",X"B1",X"48",
		X"A4",X"40",X"99",X"F8",X"04",X"8A",X"0A",X"AA",X"20",X"07",X"C9",X"B0",X"02",X"A9",X"00",X"AA",
		X"A0",X"00",X"68",X"99",X"40",X"00",X"C8",X"C0",X"0D",X"90",X"F7",X"8A",X"A0",X"02",X"A2",X"00",
		X"C9",X"01",X"60",X"A9",X"04",X"D0",X"E8",X"BD",X"1B",X"C9",X"48",X"BD",X"1A",X"C9",X"48",X"60",
		X"03",X"03",X"03",X"01",X"03",X"01",X"01",X"01",X"04",X"04",X"2D",X"C9",X"34",X"CB",X"2C",X"CB",
		X"A7",X"CA",X"2E",X"CA",X"50",X"CA",X"5A",X"CA",X"5A",X"CA",X"EF",X"C9",X"EF",X"C9",X"20",X"5F",
		X"CA",X"B0",X"37",X"A4",X"40",X"B9",X"F8",X"04",X"D0",X"38",X"A5",X"4C",X"F0",X"14",X"C9",X"49",
		X"F0",X"09",X"C9",X"48",X"D0",X"08",X"A9",X"40",X"99",X"78",X"07",X"4C",X"DB",X"C9",X"A9",X"21",
		X"38",X"60",X"A4",X"40",X"18",X"B9",X"78",X"06",X"79",X"F8",X"06",X"A0",X"00",X"91",X"4A",X"A0",
		X"07",X"B9",X"6A",X"C9",X"91",X"4A",X"88",X"D0",X"F8",X"18",X"60",X"40",X"00",X"CC",X"00",X"20",
		X"00",X"00",X"38",X"E9",X"01",X"20",X"B3",X"CD",X"B0",X"0E",X"A6",X"4C",X"F0",X"18",X"CA",X"F0",
		X"08",X"CA",X"CA",X"F0",X"11",X"A9",X"21",X"38",X"60",X"A9",X"01",X"A0",X"00",X"91",X"4A",X"A8",
		X"A9",X"00",X"91",X"4A",X"18",X"60",X"A9",X"F8",X"A0",X"00",X"91",X"4A",X"A6",X"41",X"A4",X"40",
		X"20",X"E6",X"CA",X"B0",X"C5",X"98",X"A0",X"02",X"91",X"4A",X"88",X"8A",X"91",X"4A",X"A0",X"03",
		X"A9",X"00",X"91",X"4A",X"A5",X"4C",X"F0",X"0C",X"A0",X"04",X"B9",X"C2",X"C9",X"91",X"4A",X"C8",
		X"C0",X"19",X"90",X"F6",X"18",X"60",X"10",X"43",X"4F",X"4D",X"50",X"41",X"43",X"54",X"20",X"46",
		X"4C",X"41",X"53",X"48",X"20",X"20",X"20",X"02",X"20",X"00",X"20",X"A4",X"40",X"A6",X"41",X"20",
		X"99",X"CD",X"D0",X"04",X"A9",X"28",X"38",X"60",X"20",X"2B",X"CD",X"20",X"10",X"CD",X"D0",X"04",
		X"A9",X"27",X"38",X"60",X"A0",X"01",X"84",X"42",X"88",X"BD",X"88",X"C0",X"91",X"4A",X"C8",X"BD",
		X"80",X"C0",X"91",X"4A",X"C8",X"D0",X"F2",X"E6",X"4B",X"C6",X"42",X"10",X"EC",X"C6",X"4B",X"C6",
		X"4B",X"A0",X"2E",X"A2",X"18",X"20",X"1C",X"CA",X"A0",X"14",X"A2",X"0A",X"B1",X"4A",X"48",X"C8",
		X"B1",X"4A",X"88",X"91",X"4A",X"C8",X"68",X"91",X"4A",X"C8",X"CA",X"D0",X"EF",X"18",X"60",X"20",
		X"5F",X"CA",X"B0",X"18",X"20",X"A8",X"CA",X"B0",X"13",X"A6",X"4C",X"F0",X"0F",X"CA",X"F0",X"0C",
		X"CA",X"F0",X"06",X"CA",X"F0",X"07",X"CA",X"F0",X"03",X"A9",X"21",X"38",X"60",X"A9",X"1F",X"38",
		X"60",X"B9",X"F8",X"04",X"18",X"F0",X"03",X"A9",X"11",X"38",X"60",X"A9",X"01",X"38",X"60",X"A0",
		X"02",X"B1",X"48",X"85",X"4A",X"C8",X"B1",X"48",X"85",X"4B",X"C8",X"B1",X"48",X"85",X"4C",X"18",
		X"60",X"A0",X"02",X"B1",X"48",X"85",X"44",X"C8",X"B1",X"48",X"85",X"45",X"C8",X"B1",X"48",X"85",
		X"46",X"C8",X"B1",X"48",X"85",X"47",X"A4",X"40",X"B9",X"F8",X"04",X"20",X"A8",X"CA",X"B0",X"17",
		X"A0",X"06",X"B1",X"48",X"D0",X"0E",X"A5",X"47",X"25",X"46",X"C9",X"FF",X"F0",X"06",X"A4",X"40",
		X"A6",X"41",X"18",X"60",X"A9",X"2D",X"38",X"60",X"A4",X"40",X"B9",X"F8",X"04",X"38",X"F0",X"06",
		X"38",X"E9",X"01",X"20",X"B3",X"CD",X"A9",X"11",X"60",X"90",X"03",X"4C",X"8C",X"C8",X"20",X"FB",
		X"CB",X"8A",X"45",X"43",X"29",X"70",X"F0",X"02",X"A9",X"02",X"24",X"43",X"10",X"03",X"18",X"69",
		X"01",X"20",X"B3",X"CD",X"B0",X"0E",X"A5",X"42",X"F0",X"0C",X"C9",X"01",X"F0",X"5C",X"C9",X"02",
		X"F0",X"50",X"A9",X"27",X"38",X"60",X"B9",X"78",X"07",X"0A",X"30",X"0D",X"B9",X"F8",X"04",X"18",
		X"69",X"01",X"D9",X"78",X"06",X"F0",X"15",X"D0",X"0B",X"B9",X"F8",X"04",X"18",X"69",X"01",X"D9",
		X"F8",X"06",X"F0",X"08",X"A2",X"FF",X"A0",X"FF",X"A9",X"00",X"18",X"60",X"A5",X"08",X"48",X"A5",
		X"07",X"48",X"A5",X"06",X"48",X"20",X"3B",X"CD",X"A4",X"07",X"A6",X"06",X"68",X"85",X"06",X"68",
		X"85",X"07",X"68",X"85",X"08",X"B0",X"03",X"A9",X"00",X"60",X"A9",X"27",X"60",X"20",X"71",X"CA",
		X"B0",X"FA",X"38",X"B0",X"06",X"20",X"71",X"CA",X"B0",X"F2",X"18",X"A5",X"47",X"48",X"A5",X"46",
		X"48",X"A5",X"45",X"48",X"A5",X"EF",X"48",X"08",X"20",X"BD",X"CB",X"28",X"A9",X"20",X"90",X"02",
		X"A9",X"30",X"08",X"20",X"12",X"CD",X"F0",X"60",X"28",X"A0",X"01",X"84",X"EF",X"88",X"B0",X"17",
		X"BD",X"88",X"C0",X"91",X"44",X"C8",X"BD",X"80",X"C0",X"91",X"44",X"C8",X"D0",X"F2",X"E6",X"45",
		X"C6",X"EF",X"10",X"EC",X"4C",X"A0",X"CB",X"A5",X"44",X"18",X"69",X"01",X"85",X"46",X"A5",X"45",
		X"69",X"00",X"85",X"47",X"BD",X"81",X"C0",X"B1",X"46",X"9D",X"80",X"C0",X"B1",X"44",X"9D",X"88",
		X"C0",X"C8",X"C8",X"D0",X"F2",X"E6",X"45",X"E6",X"47",X"C6",X"EF",X"10",X"EA",X"BD",X"82",X"C0",
		X"20",X"21",X"CD",X"F0",X"14",X"A9",X"00",X"C9",X"01",X"AA",X"68",X"85",X"EF",X"68",X"85",X"45",
		X"68",X"85",X"46",X"68",X"85",X"47",X"8A",X"60",X"28",X"A9",X"27",X"D0",X"EA",X"20",X"2B",X"CD",
		X"A9",X"01",X"9D",X"8A",X"C0",X"B9",X"78",X"07",X"0A",X"30",X"1A",X"A5",X"46",X"6D",X"0F",X"C8",
		X"9D",X"8B",X"C0",X"A5",X"47",X"6D",X"10",X"C8",X"9D",X"8C",X"C0",X"AD",X"11",X"C8",X"79",X"F8",
		X"04",X"9D",X"8D",X"C0",X"60",X"A5",X"46",X"6D",X"12",X"C8",X"9D",X"8B",X"C0",X"A5",X"47",X"6D",
		X"13",X"C8",X"9D",X"8C",X"C0",X"AD",X"14",X"C8",X"4C",X"DE",X"CB",X"B9",X"78",X"04",X"C9",X"A5",
		X"F0",X"49",X"AD",X"03",X"C8",X"38",X"E9",X"01",X"99",X"F8",X"07",X"AD",X"02",X"C8",X"99",X"78",
		X"05",X"AD",X"00",X"C8",X"99",X"78",X"06",X"AD",X"01",X"C8",X"99",X"F8",X"06",X"19",X"78",X"06",
		X"F0",X"24",X"BD",X"82",X"C0",X"A9",X"00",X"9D",X"80",X"C0",X"AD",X"0E",X"C8",X"30",X"14",X"A9",
		X"06",X"9D",X"86",X"C0",X"A9",X"04",X"20",X"A7",X"CD",X"A9",X"02",X"9D",X"86",X"C0",X"A9",X"7C",
		X"20",X"A7",X"CD",X"20",X"51",X"CC",X"A9",X"A5",X"99",X"78",X"04",X"A9",X"00",X"99",X"78",X"07",
		X"60",X"BD",X"82",X"C0",X"20",X"87",X"CC",X"90",X"09",X"A9",X"00",X"99",X"78",X"06",X"99",X"F8",
		X"06",X"60",X"B9",X"78",X"06",X"F0",X"0D",X"A9",X"E0",X"20",X"A9",X"CC",X"D9",X"78",X"06",X"B0",
		X"03",X"99",X"78",X"06",X"B9",X"F8",X"06",X"F0",X"0D",X"A9",X"F0",X"20",X"A9",X"CC",X"D9",X"F8",
		X"06",X"B0",X"03",X"99",X"F8",X"06",X"60",X"98",X"48",X"AC",X"0C",X"C8",X"BD",X"8F",X"C0",X"10",
		X"14",X"A9",X"0A",X"48",X"A9",X"C5",X"20",X"A7",X"CD",X"68",X"38",X"E9",X"01",X"D0",X"F4",X"88",
		X"D0",X"EA",X"38",X"B0",X"01",X"18",X"68",X"A8",X"60",X"9D",X"8E",X"C0",X"99",X"F8",X"05",X"98",
		X"48",X"AC",X"0D",X"C8",X"BD",X"8F",X"C0",X"29",X"D0",X"C9",X"50",X"F0",X"15",X"A9",X"C5",X"20",
		X"A7",X"CD",X"88",X"D0",X"EF",X"68",X"A8",X"B9",X"F8",X"05",X"49",X"10",X"9D",X"8E",X"C0",X"A9",
		X"00",X"60",X"68",X"A8",X"BD",X"8E",X"C0",X"29",X"10",X"0A",X"0A",X"99",X"78",X"07",X"A5",X"08",
		X"48",X"A5",X"07",X"48",X"A5",X"06",X"48",X"20",X"3B",X"CD",X"A9",X"00",X"B0",X"0A",X"A5",X"06",
		X"05",X"07",X"C9",X"01",X"A5",X"08",X"69",X"00",X"99",X"F8",X"05",X"68",X"85",X"06",X"68",X"85",
		X"07",X"68",X"85",X"08",X"B9",X"F8",X"05",X"60",X"BD",X"8F",X"C0",X"30",X"FB",X"29",X"08",X"60",
		X"A9",X"EC",X"48",X"BD",X"8F",X"C0",X"30",X"FB",X"A9",X"00",X"9D",X"80",X"C0",X"68",X"9D",X"8F",
		X"C0",X"BD",X"8F",X"C0",X"30",X"FB",X"29",X"09",X"C9",X"01",X"60",X"20",X"08",X"CD",X"B9",X"78",
		X"07",X"4A",X"4A",X"29",X"10",X"09",X"E0",X"9D",X"8E",X"C0",X"60",X"20",X"2B",X"CD",X"20",X"10",
		X"CD",X"D0",X"04",X"A9",X"27",X"38",X"60",X"98",X"48",X"A0",X"00",X"BD",X"88",X"C0",X"C8",X"C0",
		X"39",X"D0",X"F8",X"68",X"A8",X"B9",X"78",X"07",X"0A",X"0A",X"98",X"48",X"A0",X"00",X"90",X"02",
		X"A0",X"03",X"38",X"BD",X"88",X"C0",X"F9",X"0F",X"C8",X"85",X"06",X"BD",X"80",X"C0",X"F9",X"10",
		X"C8",X"85",X"07",X"BD",X"88",X"C0",X"F9",X"11",X"C8",X"85",X"08",X"BD",X"80",X"C0",X"E9",X"00",
		X"F0",X"08",X"A9",X"FF",X"85",X"06",X"85",X"07",X"85",X"08",X"68",X"A8",X"20",X"08",X"CD",X"F0",
		X"06",X"BD",X"88",X"C0",X"4C",X"8C",X"CD",X"18",X"60",X"B9",X"78",X"07",X"0A",X"30",X"04",X"B9",
		X"78",X"06",X"60",X"B9",X"F8",X"06",X"60",X"38",X"48",X"E9",X"01",X"D0",X"FC",X"68",X"E9",X"01",
		X"D0",X"F6",X"60",X"48",X"B9",X"78",X"05",X"D0",X"22",X"68",X"F0",X"09",X"D9",X"F8",X"07",X"D0",
		X"07",X"A9",X"00",X"F0",X"03",X"B9",X"F8",X"07",X"99",X"F8",X"04",X"38",X"F9",X"78",X"06",X"90",
		X"32",X"99",X"F8",X"04",X"D9",X"F8",X"06",X"B0",X"22",X"90",X"23",X"68",X"F0",X"09",X"D9",X"F8",
		X"07",X"D0",X"07",X"A9",X"00",X"F0",X"03",X"B9",X"F8",X"07",X"99",X"F8",X"04",X"38",X"F9",X"F8",
		X"06",X"90",X"0B",X"99",X"F8",X"04",X"D9",X"78",X"06",X"90",X"08",X"A9",X"28",X"60",X"A9",X"40",
		X"99",X"78",X"07",X"B9",X"F8",X"04",X"60",X"0A",X"0B",X"0D",X"0E",X"15",X"03",X"0E",X"0A",X"09",
		X"08",X"1C",X"2B",X"2F",X"37",X"40",X"00",X"00",X"00",X"01",X"0E",X"0E",X"02",X"0E",X"86",X"41",
		X"84",X"40",X"84",X"01",X"A9",X"00",X"8D",X"F2",X"03",X"A9",X"E0",X"8D",X"F3",X"03",X"20",X"6F",
		X"FB",X"20",X"59",X"C8",X"A6",X"41",X"A4",X"40",X"20",X"02",X"CC",X"8D",X"10",X"C0",X"A4",X"40",
		X"B9",X"78",X"05",X"85",X"87",X"B9",X"F8",X"07",X"18",X"69",X"01",X"85",X"88",X"A2",X"01",X"D0",
		X"02",X"A2",X"03",X"BD",X"00",X"C8",X"95",X"85",X"CA",X"10",X"F8",X"A9",X"03",X"85",X"82",X"A9",
		X"00",X"85",X"83",X"A2",X"04",X"BD",X"07",X"CE",X"20",X"5B",X"FB",X"BD",X"0C",X"CE",X"85",X"24",
		X"BD",X"11",X"CE",X"A8",X"20",X"61",X"CF",X"E0",X"04",X"F0",X"22",X"A0",X"13",X"20",X"61",X"CF",
		X"B5",X"85",X"DD",X"00",X"C8",X"F0",X"0A",X"E0",X"02",X"B0",X"02",X"E6",X"83",X"A0",X"3F",X"84",
		X"32",X"20",X"6D",X"CF",X"A0",X"FF",X"84",X"32",X"A9",X"A0",X"20",X"ED",X"FD",X"CA",X"10",X"C5",
		X"A4",X"40",X"A5",X"87",X"99",X"78",X"05",X"A5",X"88",X"38",X"E9",X"01",X"99",X"F8",X"07",X"A6",
		X"82",X"BD",X"07",X"CE",X"20",X"5B",X"FB",X"A9",X"16",X"85",X"24",X"D0",X"03",X"20",X"DD",X"FB",
		X"20",X"0C",X"FD",X"C9",X"9B",X"F0",X"8A",X"C9",X"88",X"D0",X"12",X"A9",X"FE",X"75",X"85",X"DD",
		X"16",X"CE",X"90",X"E9",X"DD",X"1A",X"CE",X"B0",X"E4",X"95",X"85",X"90",X"82",X"C9",X"95",X"D0",
		X"04",X"A9",X"00",X"F0",X"E8",X"C9",X"8D",X"F0",X"04",X"C9",X"8A",X"D0",X"0F",X"8A",X"18",X"69",
		X"01",X"C9",X"04",X"90",X"02",X"A9",X"00",X"85",X"82",X"4C",X"AF",X"CE",X"C9",X"8B",X"D0",X"08",
		X"C6",X"82",X"10",X"F5",X"A9",X"03",X"D0",X"EF",X"29",X"DF",X"C9",X"C2",X"D0",X"0F",X"A5",X"83",
		X"D0",X"AB",X"20",X"58",X"FC",X"AD",X"F8",X"07",X"85",X"84",X"6C",X"83",X"00",X"C9",X"D3",X"F0",
		X"0A",X"C9",X"D1",X"D0",X"D4",X"20",X"58",X"FC",X"4C",X"00",X"E0",X"A2",X"0E",X"BD",X"F0",X"CF",
		X"95",X"90",X"CA",X"10",X"F8",X"A6",X"41",X"9D",X"83",X"C0",X"A2",X"03",X"B5",X"85",X"DD",X"00",
		X"C8",X"F0",X"0E",X"E0",X"02",X"B0",X"05",X"A4",X"40",X"99",X"78",X"04",X"20",X"90",X"00",X"F0",
		X"0A",X"CA",X"10",X"E8",X"A6",X"41",X"9D",X"84",X"C0",X"D0",X"03",X"20",X"DD",X"FB",X"4C",X"5F",
		X"CE",X"B9",X"9A",X"CF",X"48",X"20",X"31",X"C8",X"C8",X"68",X"10",X"F5",X"60",X"C9",X"0A",X"90",
		X"11",X"C9",X"14",X"90",X"04",X"A9",X"3F",X"D0",X"0B",X"E9",X"09",X"48",X"A9",X"B1",X"20",X"ED",
		X"FD",X"68",X"09",X"B0",X"09",X"80",X"C9",X"E1",X"90",X"0D",X"48",X"AD",X"B3",X"FB",X"49",X"06",
		X"C9",X"01",X"68",X"90",X"02",X"29",X"DF",X"4C",X"ED",X"FD",X"43",X"46",X"46",X"41",X"20",X"36",
		X"35",X"30",X"32",X"20",X"76",X"32",X"2E",X"B0",X"53",X"6C",X"6F",X"74",X"A0",X"3A",X"A0",X"0D",
		X"0D",X"45",X"72",X"72",X"20",X"A4",X"50",X"61",X"72",X"74",X"69",X"74",X"69",X"6F",X"6E",X"73",
		X"20",X"44",X"65",X"76",X"B0",X"44",X"65",X"76",X"B1",X"42",X"6F",X"6F",X"74",X"20",X"44",X"65",
		X"F6",X"50",X"61",X"72",X"74",X"69",X"74",X"69",X"6F",X"EE",X"42",X"29",X"4F",X"4F",X"54",X"20",
		X"53",X"29",X"41",X"56",X"45",X"20",X"51",X"29",X"55",X"49",X"D4",X"77",X"77",X"77",X"77",X"FF",
		X"9D",X"00",X"C8",X"A0",X"00",X"88",X"F0",X"05",X"DD",X"00",X"C8",X"D0",X"F8",X"98",X"60",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
