library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ssc_rom is
port (
	clk  : in  std_logic;
	addr : in  unsigned(10 downto 0);
	data : out unsigned(7 downto 0)
);
end entity;

architecture prom of ssc_rom is
	type rom is array(0 to  2047) of unsigned(7 downto 0);
	signal rom_data: rom := (
		X"20",X"9B",X"C9",X"A9",X"16",X"48",X"A9",X"00",X"9D",X"B8",X"04",X"9D",X"B8",X"03",X"9D",X"38",
		X"04",X"9D",X"B8",X"05",X"9D",X"38",X"06",X"9D",X"B8",X"06",X"B9",X"82",X"C0",X"85",X"2B",X"4A",
		X"4A",X"90",X"04",X"68",X"29",X"FE",X"48",X"B8",X"B9",X"81",X"C0",X"4A",X"B0",X"07",X"4A",X"B0",
		X"0E",X"A9",X"01",X"D0",X"3D",X"4A",X"A9",X"03",X"B0",X"02",X"A9",X"80",X"9D",X"B8",X"04",X"2C",
		X"58",X"FF",X"A5",X"2B",X"29",X"20",X"49",X"20",X"9D",X"B8",X"03",X"70",X"0A",X"20",X"9B",X"C8",
		X"AE",X"F8",X"07",X"9D",X"B8",X"05",X"60",X"A5",X"2B",X"4A",X"4A",X"29",X"03",X"A8",X"F0",X"04",
		X"68",X"29",X"7F",X"48",X"B9",X"A6",X"C9",X"9D",X"38",X"06",X"A4",X"26",X"68",X"29",X"95",X"48",
		X"A9",X"09",X"9D",X"38",X"05",X"68",X"9D",X"38",X"07",X"A5",X"2B",X"48",X"29",X"A0",X"50",X"02",
		X"29",X"80",X"20",X"A1",X"CD",X"20",X"81",X"CD",X"68",X"29",X"0C",X"50",X"02",X"A9",X"00",X"0A",
		X"0A",X"0A",X"09",X"0B",X"99",X"8A",X"C0",X"B9",X"88",X"C0",X"60",X"20",X"9B",X"C9",X"20",X"AA",
		X"C8",X"29",X"7F",X"AC",X"F8",X"07",X"BE",X"B8",X"05",X"60",X"20",X"FF",X"CA",X"B0",X"05",X"20",
		X"2C",X"CC",X"90",X"F6",X"60",X"20",X"1E",X"CA",X"68",X"A8",X"68",X"AA",X"A5",X"27",X"60",X"F0",
		X"29",X"BD",X"B8",X"06",X"10",X"05",X"5E",X"B8",X"06",X"D0",X"24",X"20",X"3E",X"CC",X"90",X"1A",
		X"BD",X"B8",X"03",X"29",X"C0",X"F0",X"0E",X"A5",X"27",X"C9",X"E0",X"90",X"08",X"BD",X"B8",X"04",
		X"09",X"40",X"9D",X"B8",X"04",X"28",X"F0",X"D0",X"D0",X"CB",X"20",X"FF",X"CA",X"90",X"DC",X"20",
		X"11",X"CC",X"28",X"08",X"F0",X"DA",X"20",X"D1",X"C9",X"4C",X"D0",X"C8",X"20",X"1A",X"CB",X"B0",
		X"B7",X"A5",X"27",X"48",X"BD",X"38",X"07",X"29",X"C0",X"D0",X"16",X"A5",X"24",X"F0",X"42",X"C9",
		X"08",X"F0",X"04",X"C9",X"10",X"D0",X"0A",X"09",X"F0",X"3D",X"B8",X"06",X"18",X"65",X"24",X"85",
		X"24",X"BD",X"B8",X"06",X"C5",X"24",X"F0",X"29",X"A9",X"A0",X"90",X"08",X"BD",X"38",X"07",X"0A",
		X"10",X"1F",X"A9",X"88",X"85",X"27",X"2C",X"58",X"FF",X"08",X"70",X"0C",X"EA",X"2C",X"58",X"FF",
		X"50",X"B8",X"AE",X"F8",X"07",X"4C",X"EF",X"C9",X"20",X"B5",X"C9",X"20",X"6B",X"CB",X"4C",X"68",
		X"C9",X"68",X"B8",X"08",X"85",X"27",X"48",X"20",X"68",X"CB",X"20",X"B5",X"C9",X"68",X"49",X"8D",
		X"0A",X"D0",X"05",X"9D",X"B8",X"06",X"85",X"24",X"BD",X"B8",X"04",X"10",X"0D",X"BD",X"38",X"06",
		X"F0",X"08",X"18",X"FD",X"B8",X"06",X"A9",X"8D",X"90",X"DA",X"28",X"70",X"A4",X"BD",X"38",X"07",
		X"30",X"16",X"BC",X"B8",X"06",X"0A",X"30",X"0E",X"98",X"A0",X"00",X"38",X"FD",X"38",X"06",X"C9",
		X"F8",X"90",X"03",X"69",X"27",X"A8",X"84",X"24",X"4C",X"B8",X"C8",X"8E",X"F8",X"07",X"84",X"26",
		X"A9",X"00",X"9D",X"B8",X"05",X"60",X"29",X"48",X"50",X"84",X"85",X"27",X"20",X"9B",X"C9",X"20",
		X"63",X"CB",X"4C",X"A3",X"C8",X"A5",X"27",X"49",X"08",X"0A",X"F0",X"04",X"49",X"EE",X"D0",X"09",
		X"DE",X"B8",X"06",X"10",X"03",X"9D",X"B8",X"06",X"60",X"C9",X"C0",X"B0",X"FB",X"FE",X"B8",X"06",
		X"60",X"BD",X"38",X"07",X"29",X"08",X"F0",X"16",X"BD",X"B8",X"04",X"A4",X"27",X"C0",X"94",X"D0",
		X"04",X"09",X"80",X"D0",X"06",X"C0",X"92",X"D0",X"05",X"29",X"7F",X"9D",X"B8",X"04",X"60",X"8A",
		X"0A",X"0A",X"0A",X"0A",X"85",X"26",X"A9",X"00",X"9D",X"B8",X"05",X"70",X"0F",X"A0",X"00",X"B1",
		X"3C",X"85",X"27",X"20",X"02",X"CC",X"20",X"BA",X"FC",X"90",X"F2",X"60",X"20",X"D2",X"CA",X"90",
		X"FB",X"B9",X"88",X"C0",X"A0",X"00",X"91",X"3C",X"20",X"BA",X"FC",X"90",X"EF",X"60",X"BD",X"B8",
		X"04",X"10",X"31",X"A9",X"02",X"48",X"A9",X"7F",X"20",X"E2",X"CD",X"A4",X"24",X"B1",X"28",X"85",
		X"27",X"A9",X"07",X"25",X"4F",X"D0",X"10",X"A4",X"24",X"A9",X"DF",X"D1",X"28",X"D0",X"02",X"A5",
		X"27",X"91",X"28",X"E6",X"4F",X"E6",X"4F",X"BD",X"B8",X"04",X"30",X"09",X"20",X"11",X"CC",X"68",
		X"A9",X"8D",X"85",X"27",X"60",X"20",X"FF",X"CA",X"90",X"0C",X"20",X"11",X"CC",X"20",X"D1",X"C9",
		X"20",X"A3",X"CC",X"4C",X"2B",X"CA",X"20",X"3E",X"CC",X"90",X"C6",X"70",X"BE",X"BD",X"38",X"07",
		X"0A",X"10",X"22",X"68",X"A8",X"A5",X"27",X"C0",X"01",X"F0",X"20",X"B0",X"34",X"C9",X"9B",X"D0",
		X"06",X"C8",X"98",X"48",X"4C",X"2B",X"CA",X"C9",X"C1",X"90",X"08",X"C9",X"DB",X"B0",X"04",X"09",
		X"20",X"85",X"27",X"98",X"48",X"20",X"68",X"CB",X"4C",X"2B",X"CA",X"C9",X"9B",X"F0",X"E2",X"C9",
		X"B0",X"90",X"0A",X"C9",X"BB",X"B0",X"06",X"A8",X"B9",X"09",X"CA",X"85",X"27",X"A0",X"00",X"F0",
		X"E2",X"C9",X"9B",X"D0",X"DE",X"A0",X"00",X"F0",X"C9",X"9B",X"9C",X"9F",X"DB",X"DC",X"DF",X"FB",
		X"FC",X"FD",X"FE",X"FF",X"A2",X"CA",X"CA",X"D0",X"FD",X"38",X"E9",X"01",X"D0",X"F6",X"AE",X"F8",
		X"07",X"60",X"A4",X"26",X"B9",X"89",X"C0",X"48",X"29",X"20",X"4A",X"4A",X"85",X"35",X"68",X"29",
		X"0F",X"C9",X"08",X"90",X"04",X"29",X"07",X"B0",X"02",X"A5",X"35",X"05",X"35",X"F0",X"05",X"09",
		X"20",X"9D",X"B8",X"05",X"60",X"A4",X"26",X"B9",X"89",X"C0",X"29",X"70",X"C9",X"10",X"60",X"20",
		X"D2",X"CA",X"90",X"15",X"B9",X"88",X"C0",X"09",X"80",X"C9",X"8A",X"D0",X"09",X"A8",X"BD",X"38",
		X"07",X"29",X"20",X"D0",X"03",X"98",X"38",X"60",X"18",X"60",X"A4",X"26",X"B9",X"81",X"C0",X"4A",
		X"B0",X"36",X"BD",X"B8",X"04",X"29",X"07",X"F0",X"05",X"20",X"FC",X"CD",X"38",X"60",X"A5",X"27",
		X"29",X"7F",X"DD",X"38",X"05",X"D0",X"05",X"FE",X"B8",X"04",X"38",X"60",X"BD",X"38",X"07",X"29",
		X"08",X"F0",X"15",X"20",X"FF",X"CA",X"90",X"10",X"C9",X"93",X"F0",X"0E",X"48",X"BD",X"38",X"07",
		X"4A",X"4A",X"68",X"90",X"04",X"9D",X"B8",X"06",X"18",X"60",X"20",X"AA",X"C8",X"C9",X"91",X"D0",
		X"F9",X"18",X"60",X"20",X"1A",X"CB",X"B0",X"F1",X"20",X"9E",X"CC",X"A4",X"26",X"B9",X"81",X"C0",
		X"4A",X"90",X"4E",X"4A",X"90",X"4B",X"A5",X"27",X"48",X"BD",X"38",X"04",X"C9",X"67",X"90",X"10",
		X"C9",X"6C",X"B0",X"22",X"C9",X"6B",X"68",X"48",X"49",X"9B",X"29",X"7F",X"D0",X"18",X"B0",X"19",
		X"BD",X"B8",X"04",X"29",X"1F",X"09",X"80",X"85",X"27",X"20",X"02",X"CC",X"20",X"AA",X"C8",X"49",
		X"86",X"D0",X"ED",X"9D",X"38",X"04",X"DE",X"38",X"04",X"68",X"85",X"27",X"49",X"8D",X"0A",X"D0",
		X"0A",X"BD",X"B8",X"03",X"29",X"30",X"F0",X"03",X"9D",X"38",X"04",X"20",X"02",X"CC",X"4C",X"EA",
		X"CB",X"20",X"02",X"CC",X"0A",X"A8",X"BD",X"B8",X"03",X"C0",X"18",X"F0",X"0C",X"4A",X"4A",X"C0",
		X"14",X"F0",X"06",X"4A",X"4A",X"C0",X"1A",X"D0",X"25",X"29",X"03",X"F0",X"0D",X"A8",X"B9",X"FE",
		X"CB",X"A8",X"A9",X"20",X"20",X"C4",X"CA",X"88",X"D0",X"F8",X"A5",X"27",X"0A",X"C9",X"1A",X"D0",
		X"0D",X"BD",X"38",X"07",X"6A",X"90",X"07",X"A9",X"8A",X"85",X"27",X"4C",X"6B",X"CB",X"60",X"01",
		X"08",X"40",X"20",X"F5",X"CA",X"D0",X"FB",X"98",X"09",X"89",X"A8",X"A5",X"27",X"99",X"FF",X"BF",
		X"60",X"48",X"A4",X"24",X"A5",X"27",X"91",X"28",X"68",X"C9",X"95",X"D0",X"0C",X"A5",X"27",X"C9",
		X"20",X"B0",X"06",X"20",X"DF",X"CC",X"59",X"DB",X"CC",X"85",X"27",X"60",X"18",X"BD",X"38",X"07",
		X"29",X"04",X"F0",X"09",X"AD",X"00",X"C0",X"10",X"04",X"8D",X"10",X"C0",X"38",X"60",X"E6",X"4E",
		X"D0",X"02",X"E6",X"4F",X"20",X"2C",X"CC",X"B8",X"90",X"F3",X"20",X"11",X"CC",X"29",X"7F",X"DD",
		X"38",X"05",X"D0",X"3D",X"A4",X"26",X"B9",X"81",X"C0",X"4A",X"B0",X"35",X"A0",X"0A",X"B9",X"93",
		X"CC",X"85",X"27",X"98",X"48",X"20",X"A3",X"CC",X"68",X"A8",X"88",X"10",X"F1",X"A9",X"01",X"20",
		X"7B",X"CE",X"20",X"34",X"CC",X"10",X"FB",X"C9",X"88",X"F0",X"E1",X"85",X"27",X"20",X"A3",X"CC",
		X"20",X"1A",X"CB",X"BD",X"B8",X"04",X"29",X"07",X"D0",X"E8",X"A9",X"8D",X"85",X"27",X"2C",X"58",
		X"FF",X"38",X"60",X"BA",X"C3",X"D3",X"D3",X"A0",X"C5",X"CC",X"D0",X"D0",X"C1",X"8D",X"BD",X"38",
		X"07",X"10",X"13",X"BD",X"38",X"07",X"29",X"02",X"F0",X"0D",X"BD",X"B8",X"04",X"29",X"38",X"F0",
		X"06",X"8A",X"48",X"A9",X"AF",X"48",X"60",X"20",X"DF",X"CC",X"09",X"80",X"C9",X"E0",X"90",X"06",
		X"59",X"D3",X"CC",X"4C",X"F6",X"FD",X"C9",X"C1",X"90",X"F9",X"C9",X"DB",X"B0",X"F5",X"59",X"D7",
		X"CC",X"90",X"F0",X"20",X"00",X"E0",X"20",X"00",X"00",X"00",X"C0",X"00",X"00",X"E0",X"C0",X"BD",
		X"B8",X"03",X"2A",X"2A",X"2A",X"29",X"03",X"A8",X"A5",X"27",X"60",X"42",X"67",X"C0",X"54",X"47",
		X"A6",X"43",X"87",X"A6",X"51",X"47",X"B8",X"52",X"C7",X"AC",X"5A",X"E7",X"F3",X"49",X"90",X"D3",
		X"4B",X"90",X"DF",X"45",X"43",X"80",X"46",X"E3",X"04",X"4C",X"E3",X"01",X"58",X"E3",X"08",X"54",
		X"83",X"40",X"53",X"43",X"40",X"4D",X"E3",X"20",X"00",X"42",X"F6",X"7C",X"50",X"F6",X"9A",X"44",
		X"F6",X"9B",X"46",X"F6",X"46",X"4C",X"F6",X"40",X"43",X"F6",X"3A",X"54",X"D6",X"34",X"4E",X"90",
		X"E8",X"53",X"56",X"60",X"00",X"A9",X"3F",X"A0",X"07",X"D0",X"10",X"A9",X"CF",X"A0",X"05",X"D0",
		X"0A",X"A9",X"F3",X"A0",X"03",X"D0",X"04",X"A9",X"FC",X"A0",X"01",X"3D",X"B8",X"03",X"85",X"2A",
		X"BD",X"38",X"04",X"29",X"03",X"18",X"6A",X"2A",X"88",X"D0",X"FC",X"05",X"2A",X"9D",X"B8",X"03",
		X"60",X"29",X"07",X"0A",X"0A",X"0A",X"85",X"2A",X"0A",X"C5",X"26",X"F0",X"0F",X"BD",X"B8",X"04",
		X"29",X"C7",X"05",X"2A",X"9D",X"B8",X"04",X"A9",X"00",X"9D",X"38",X"06",X"60",X"29",X"0F",X"D0",
		X"07",X"B9",X"81",X"C0",X"4A",X"4A",X"4A",X"4A",X"09",X"10",X"85",X"2A",X"A9",X"E0",X"85",X"2B",
		X"B9",X"8B",X"C0",X"25",X"2B",X"05",X"2A",X"99",X"8B",X"C0",X"60",X"88",X"0A",X"0A",X"0A",X"0A",
		X"0A",X"85",X"2A",X"A9",X"1F",X"D0",X"E7",X"1E",X"B8",X"04",X"38",X"B0",X"10",X"99",X"89",X"C0",
		X"20",X"93",X"FE",X"20",X"89",X"FE",X"AE",X"F8",X"07",X"1E",X"B8",X"04",X"18",X"7E",X"B8",X"04",
		X"60",X"B9",X"8A",X"C0",X"48",X"09",X"0C",X"99",X"8A",X"C0",X"A9",X"E9",X"20",X"C4",X"CA",X"68",
		X"99",X"8A",X"C0",X"60",X"A9",X"28",X"9D",X"38",X"06",X"A9",X"80",X"1D",X"38",X"07",X"D0",X"05",
		X"A9",X"FE",X"3D",X"38",X"07",X"9D",X"38",X"07",X"60",X"C9",X"28",X"90",X"0E",X"9D",X"38",X"06",
		X"A9",X"3F",X"D0",X"EE",X"1E",X"38",X"05",X"38",X"7E",X"38",X"05",X"60",X"A8",X"A5",X"27",X"29",
		X"7F",X"C9",X"20",X"D0",X"09",X"C0",X"03",X"F0",X"01",X"60",X"A9",X"04",X"D0",X"6D",X"C9",X"0D",
		X"D0",X"12",X"20",X"79",X"CE",X"C0",X"07",X"F0",X"01",X"60",X"A9",X"CD",X"48",X"BD",X"38",X"04",
		X"48",X"A4",X"26",X"60",X"85",X"35",X"A9",X"CE",X"48",X"B9",X"30",X"CE",X"48",X"A5",X"35",X"60",
		X"A7",X"37",X"61",X"89",X"8A",X"A7",X"89",X"89",X"DD",X"38",X"05",X"D0",X"06",X"DE",X"B8",X"04",
		X"4C",X"02",X"CC",X"C9",X"30",X"90",X"0D",X"C9",X"3A",X"B0",X"09",X"29",X"0F",X"9D",X"38",X"04",
		X"A9",X"02",X"D0",X"27",X"C9",X"20",X"B0",X"06",X"9D",X"38",X"05",X"4C",X"79",X"CE",X"A0",X"00",
		X"F0",X"4D",X"49",X"30",X"C9",X"0A",X"B0",X"0D",X"A0",X"0A",X"7D",X"38",X"04",X"88",X"D0",X"FA",
		X"9D",X"38",X"04",X"F0",X"15",X"A0",X"2E",X"D0",X"36",X"A9",X"00",X"85",X"2A",X"AE",X"F8",X"07",
		X"BD",X"B8",X"04",X"29",X"F8",X"05",X"2A",X"9D",X"B8",X"04",X"60",X"A8",X"BD",X"38",X"04",X"C0",
		X"44",X"F0",X"09",X"C0",X"45",X"D0",X"11",X"1D",X"38",X"07",X"D0",X"05",X"49",X"FF",X"3D",X"38",
		X"07",X"9D",X"38",X"07",X"A9",X"06",X"D0",X"D3",X"A9",X"20",X"9D",X"B8",X"05",X"D0",X"F5",X"B9",
		X"EB",X"CC",X"F0",X"F4",X"C5",X"35",X"F0",X"05",X"C8",X"C8",X"C8",X"D0",X"F2",X"C8",X"B9",X"EB",
		X"CC",X"85",X"2A",X"29",X"20",X"D0",X"07",X"BD",X"38",X"07",X"29",X"10",X"D0",X"EB",X"BD",X"38",
		X"07",X"4A",X"4A",X"24",X"2A",X"B0",X"04",X"10",X"E0",X"30",X"02",X"50",X"DC",X"A5",X"2A",X"48",
		X"29",X"07",X"20",X"7B",X"CE",X"C8",X"68",X"29",X"10",X"D0",X"07",X"B9",X"EB",X"CC",X"9D",X"38",
		X"04",X"60",X"A9",X"CD",X"48",X"B9",X"EB",X"CC",X"48",X"A4",X"26",X"BD",X"38",X"04",X"60",X"C2",
		X"2C",X"58",X"FF",X"70",X"0C",X"38",X"90",X"18",X"B8",X"50",X"06",X"01",X"31",X"8E",X"94",X"97",
		X"9A",X"85",X"27",X"86",X"35",X"8A",X"48",X"98",X"48",X"08",X"78",X"8D",X"FF",X"CF",X"20",X"58",
		X"FF",X"BA",X"BD",X"00",X"01",X"8D",X"F8",X"07",X"AA",X"0A",X"0A",X"0A",X"0A",X"85",X"26",X"A8",
		X"28",X"50",X"29",X"1E",X"38",X"05",X"5E",X"38",X"05",X"B9",X"8A",X"C0",X"29",X"1F",X"D0",X"05",
		X"A9",X"EF",X"20",X"05",X"C8",X"E4",X"37",X"D0",X"0B",X"A9",X"07",X"C5",X"36",X"F0",X"05",X"85",
		X"36",X"18",X"90",X"08",X"E4",X"39",X"D0",X"F9",X"A9",X"05",X"85",X"38",X"BD",X"38",X"07",X"29",
		X"02",X"08",X"90",X"03",X"4C",X"BF",X"C8",X"BD",X"B8",X"04",X"48",X"0A",X"10",X"0E",X"A6",X"35",
		X"A5",X"27",X"09",X"20",X"9D",X"00",X"02",X"85",X"27",X"AE",X"F8",X"07",X"68",X"29",X"BF",X"9D",
		X"B8",X"04",X"28",X"F0",X"06",X"20",X"63",X"CB",X"4C",X"B5",X"C8",X"4C",X"FC",X"C8",X"20",X"00",
		X"C8",X"A2",X"00",X"60",X"4C",X"9B",X"C8",X"4C",X"AA",X"C9",X"4A",X"20",X"9B",X"C9",X"B0",X"08",
		X"20",X"F5",X"CA",X"F0",X"06",X"18",X"90",X"03",X"20",X"D2",X"CA",X"BD",X"B8",X"05",X"AA",X"60",
		X"A2",X"03",X"B5",X"36",X"48",X"CA",X"10",X"FA",X"AE",X"F8",X"07",X"BD",X"38",X"06",X"85",X"36",
		X"BD",X"B8",X"04",X"29",X"38",X"4A",X"4A",X"4A",X"09",X"C0",X"85",X"37",X"8A",X"48",X"A5",X"27",
		X"48",X"09",X"80",X"20",X"ED",X"FD",X"68",X"85",X"27",X"68",X"8D",X"F8",X"07",X"AA",X"0A",X"0A",
		X"0A",X"0A",X"85",X"26",X"8D",X"FF",X"CF",X"A5",X"36",X"9D",X"38",X"06",X"A2",X"00",X"68",X"95",
		X"36",X"E8",X"E0",X"04",X"90",X"F8",X"AE",X"F8",X"07",X"60",X"C1",X"D0",X"D0",X"CC",X"C5",X"08");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(addr));
	end if;
end process;
end architecture;
